*DL4736A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*6.8V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4736A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  6.261
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=123P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=149U RS=1.05 N=3.5)
.ENDS