*ZMU120 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*120V 1W Si Zener pkg:DL-41 1,2
.SUBCKT ZMU120   1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  118.4
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=22.9P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.24M RS=99 N=45)
.ENDS