*DL5241B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*11V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5241B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  10.31
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=58.2P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.94M RS=6.6 N=12)
.ENDS