*
.SUBCKT 1PS74SB23 1 2
* The Resistor R1 does not reflect
* a physical device.  Instead it
* improves modeling in the reverse
* mode of operation.
R1 1 2 2.56E+05
D1 1 2 D1PS74SB23
.MODEL D1PS74SB23 D
+(
+ IS = 6.984E-06
+ N = 1.023
+ BV = 30
+ IBV = 0.0002402
+ RS = 0.1574
+ CJO = 3.075E-10
+ VJ = 0.6615
+ M = 0.6098
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*