*SI4948EY  MCE  5-28-97
* jjt 4/4/2002: changed VTO to -1V to match  S-57253�Rev. D, 24-Feb-98 datasheet
*60V 3A 0.112ohm Dual Power MOSFET pkg:SMD8A (A:8,2,1)(B:6,4,3)
.SUBCKT SI4948EY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  52.2M
RS  40  3  3.8M
RG  20  2  48.4
CGS  2  3  1.07N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  435P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=125K THETA=80M ETA=2M VTO=-1 KP=25.2)
.MODEL DCGD D (CJO=435P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=12.9N N=1.5 RS=16.1M BV=60 CJO=417P VJ=0.8 M=0.42 TT=60N)
.MODEL DLIM D (IS=100U)
.ENDS 