*DL4738A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*8.2V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4738A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  7.658
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=92.8P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=185U RS=1.35 N=3.8)
.ENDS