*Si6956DQ Siliconix 13-Oct-96
*N-Channel DMOS Subcircuit Model
.SUBCKT Si6956DQ 4 1 2 2
M1 3 1 2 2 NMOS W=283290U L=0.5U
R1 4 3 RTEMP 32.5M
CGS 1 2 75PF
CGD 1 6 500PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=50N RS=13M RD=0 LD=0
+ NSUB=1.965E+17 UO=420 VMAX=0 ETA=1.1M XJ=500N THETA=200M
+ KAPPA=0.05 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0 IS=0)
.MODEL DMIN D(CJO=480P VJ=0.3 M=0.55 FC=0.5)
.MODEL DMAX D(CJO=240P VJ=0.9 M=0.4 FC=0.5 IS=1E-23)
.MODEL DBODY D(CJO=380P VJ=0.35 M=0.3 FC=0.5 N=1 IS=1E-10
+ TT=14N BV=30)
.MODEL RTEMP R(TC1=8M TC2=0)
.ENDS 