*SI6954DQ  MCE  5-27-97
*30V 4A 0.091ohm Dual Power MOSFET pkg:SMD8B (A:1,4,3)(B:8,5,6)
.SUBCKT SI6954DQ 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  42.2M
RS  40  3  3.28M
RG  20  2  38.5
CGS  2  3  530P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  275P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=1 KP=24.4)
.MODEL DCGD D (CJO=275P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=16.2N N=1.5 RS=5.13M BV=30 CJO=525P VJ=0.8 M=0.42 TT=48N)
.MODEL DLIM D (IS=100U)
.ENDS 