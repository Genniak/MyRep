*DL5248B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*18V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5248B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  17.46
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=41.4P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=32.6U RS=5.7 N=3.6)
.ENDS