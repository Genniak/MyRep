*ZY22 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*22V 2W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZY22     1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  21.35
.MODEL DF D (IS=10N RS=21M N=1.7 CJO=101P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.72M RS=4.5 N=10)
.ENDS