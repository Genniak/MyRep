*1N5245B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*15V 500mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5245B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  14.46
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=78.3P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=44.5U RS=4.8 N=3.7)
.ENDS