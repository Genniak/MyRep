*SI9802DY  MCE  5-27-97
*20V 4A 0.049ohm Dual Reduced Qg Power MOSFET pkg:SMD8B (A:8,2,1)(B:6,4,3)
.SUBCKT SI9802DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  22.3M
RS  40  3  2.23M
RG  20  2  33.3
CGS  2  3  490P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  476P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=41.7K THETA=80M ETA=2M VTO=0.6 KP=73.1)
.MODEL DCGD D (CJO=476P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=204N N=1.5 RS=16.2M BV=20 CJO=993P VJ=0.8 M=0.42 TT=60N)
.MODEL DLIM D (IS=100U)
.ENDS 