*DZ23C4V7 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*4.7V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C4V7 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C4V7
XB 3 2 DDZ23C4V7
.ENDS DZ23C4V7


.SUBCKT DDZ23C4V7 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  4.037
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=74.9P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=838U RS=24 N=11)
.ENDS DDZ23C4V7