*Si6433DQ Siliconix 12-Sep-94
*P-Channel DMOS Subcircuit Model
.SUBCKT Si6433DQ 4 1 2 2
M1 3 1 2 2 PMOS W=901600U L=0.5U
R1 4 3 RTEMP 18M
CGS 1 2 170PF
CGD 1 6 1450PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=17.5N RS=5.5M RD=0 LD=0 NFS=1E+12
+ NSUB=1E+16 VTO=-1.495 UO=200 VMAX=430K ETA=710U XJ=500N
+ KAPPA=1M THETA=0 TPG=-1 IS=0 KP=10.9U)
.MODEL DMIN D(CJO=3100P VJ=0.1 M=0.51 FC=0.5 IS=12E-12)
.MODEL DMAX D(CJO=3000P VJ=0.1 M=0.45 FC=0.5 IS=0.8E-20)
.MODEL DBODY D(CJO=1200P VJ=0.2 M=0.3 FC=0.5 N=1 IS=1E-10
+ TT=1.4E-7 BV=15)
.MODEL RTEMP R(TC1=3M TC2=1U)
.ENDS Si6433DQ