*Si9933DY Siliconix 16-May-95
*P-Channel DMOS Subcircuit Model
.SUBCKT Si9933DY 4 1 2 2
M1 3 1 2 2 PMOS W=547200U L=0.5U
R1 4 3 RTEMP 58M
CGS 1 2 140PF
CGD 1 6 2300PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=30N RS=20M RD=0 LD=0 NFS=1E+10
+ NSUB=1E+16 VTO=-1.7 UO=218 VMAX=400K ETA=7M XJ=800N THETA=0.1
+ KAPPA=5M CGBO=0 TPG=-1 DELTA=0.1 CGSO=0 CGDO=0 IS=0 PHI=0.18)
.MODEL DMIN D(CJO=960P VJ=0.5 M=0.9 FC=0.5 IS=1E-21)
.MODEL DMAX D(CJO=1200P VJ=0.5 M=0.5 FC=0.5 IS=1E-14 TT=10N)
.MODEL DBODY D(CJO=540P VJ=0.504 M=0.3 FC=0.5 N=1 IS=1E-12
+ TT=80N BV=16)
.MODEL RTEMP R(TC1=3M TC2=10U)
.ENDS Si9933DY