*Si6426DQ Siliconix 18-Jul-95
*N-Channel DMOS Subcircuit Model
.SUBCKT Si6426DQ 4 1 2 2
M1 3 1 2 2 NMOS W=832624U L=0.5U
R1 4 3 RTEMP 18M
CGS 1 2 905PF
CGD 1 6 2950PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=17.5N RS=500U RD=0 LD=0
+ NSUB=3.365E+17 UO=800 VMAX=2MEG ETA=300U XJ=500N
+ KAPPA=0.55 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=60.3U NFS=0.8E+12)
.MODEL DMIN D(CJO=2600P VJ=0.06 M=0.55 FC=0.5 IS=1E-20)
.MODEL DMAX D(CJO=2400P VJ=0.6 M=0.5 FC=0.5 IS=1E-16)
.MODEL DBODY D(CJO=1200P VJ=0.1 M=0.26 FC=0.5 N=1 IS=1E-15
+ TT=14N BV=40)
.MODEL RTEMP R(TC1=3.6M TC2=12U)
.ENDS 