*DZ23C20 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*20V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C20 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C20
XB 3 2 DDZ23C20
.ENDS DZ23C20


.SUBCKT DDZ23C20  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  19.4
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=31.6P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=372U RS=16.5 N=7.4)
.ENDS DDZ23C20