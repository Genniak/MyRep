*SI4425DY  MCE  5-28-97
*30V 11A 0.013ohm Power MOSFET pkg:SMD8A 5,4,1
.SUBCKT SI4425DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  5.17M
RS  40  3  1.32M
RG  20  2  13.6
CGS  2  3  4.4N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  4.13N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=-1 KP=241)
.MODEL DCGD D (CJO=4.13N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=45.7N N=1.5 RS=33.2M BV=30 CJO=1.51N VJ=0.8 M=0.42 TT=49N)
.MODEL DLIM D (IS=100U)
.ENDS 