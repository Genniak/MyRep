*1N5354B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*17V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5354B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  16.45
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=70.9P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.18M RS=0.75 N=4.7)
.ENDS