*DL4735A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*6.2V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4735A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  5.676
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=141P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=6.76U RS=0.6 N=2.2)
.ENDS