*1N4757A MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*51V 1000mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N4757A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  50.29
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=33.6P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.11M RS=28.5 N=13)
.ENDS