*1N4759A MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*62V 1000mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N4759A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  61.27
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=30.3P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=959U RS=37.5 N=14)
.ENDS