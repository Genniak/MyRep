*1N5374B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*75V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5374B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  74
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=27.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=9.04M RS=13.5 N=24)
.ENDS