*DL4741A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*11V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4741A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  10.44
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=101P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=474U RS=2.4 N=5)
.ENDS