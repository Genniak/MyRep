*SI6459DQ  MCE  5-28-97
* jjt 4/4/2002: changed sign of VTO to match S-49520�Rev. C, 18-Dec-96 datasheet.
*60V 3A 0.112ohm Power MOSFET pkg:SMD8B 1,4,6
.SUBCKT SI6459DQ 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  52.2M
RS  40  3  3.8M
RG  20  2  57.7
CGS  2  3  1E+03P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  725P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=125K THETA=80M ETA=2M VTO=-1 KP=30.1)
.MODEL DCGD D (CJO=725P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=10.8N N=1.5 RS=19.2M BV=60 CJO=463P VJ=0.8 M=0.42 TT=60N)
.MODEL DLIM D (IS=100U)
.ENDS 