*
.SUBCKT BAT120C 1 3 4
* The resistors do not reflect
* physical devices.  Instead they
* improve modeling in the reverse
* mode of operation.
R1 1 4 2.56E+05
D1 1 4 BAT120C
R2 3 4 2.56E+05
D2 3 4 BAT120C

.MODEL BAT120C D
+(
+ IS = 6.984E-06
+ N = 1.023
+ BV = 30
+ IBV = 0.0002402
+ RS = 0.1574
+ CJO = 3.075E-10
+ VJ = 0.6615
+ M = 0.6098
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*