*
* D1PS88SB48
* The resistors do not reflect
* physical devices.  Instead
* they improve modeling in the
* reverse mode of operation.
*
.SUBCKT D1PS88SB48 1 2 3
R1 1 3 8.961E+08
D1 1 3 D1PS88SB48
R2 2 3 8.961E+08
D2 2 3 D1PS88SB48
.MODEL D1PS88SB48 D
+(
+ IS = 9.649E-09
+ N = 1.013
+ BV = 1000
+ IBV = 0.001
+ RS = 4.999
+ CJO = 3.928E-12
+ VJ = 0.2057
+ M = 0.3426
+ FC = 4.441E-16
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS