*DL5237B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*8.2V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5237B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  7.664
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=46.4P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=52U RS=1.8 N=3.2)
.ENDS