*DZ23C47 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*47V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C47 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C47
XB 3 2 DDZ23C47
.ENDS DZ23C47


.SUBCKT DDZ23C47  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  46.37
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=22.1P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=245U RS=51 N=9.2)
.ENDS DDZ23C47