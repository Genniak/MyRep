*SUP75N06-08 Siliconix 07-Feb-95
*N-Channel DMOS Subcircuit Model
.SUBCKT SUP75N06-08 4 1 2 2
M1 3 1 2 2 NMOS W=8310000U L=0.5U
R1 4 3 RTEMP 4.9M
CGS 1 2 3354PF
CGD 1 6 2400PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=80N RS=1.45M RD=0 LD=0
+ NSUB=1.55E+17 UO=380 VMAX=0 ETA=0.1M XJ=500N THETA=20M
+ KAPPA=8M CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0 IS=0 NFS=3E+10)
.MODEL DMIN D(CJO=4000P VJ=0.1 M=0.53 FC=0.5 IS=1E-20 TT=10N)
.MODEL DMAX D(CJO=4000P VJ=0.9 M=0.79 FC=0.5 IS=1E-22 TT=1N)
.MODEL DBODY D(CJO=3500P VJ=0.22 M=0.36 FC=0.5 N=1 IS=1E-15
+ TT=14N BV=68)
.MODEL RTEMP R(TC1=7.55M TC2=12U)
.ENDS 