*DL4744A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*15V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4744A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  14.42
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=78.3P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=845U RS=4.2 N=6.4)
.ENDS