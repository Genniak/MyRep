*
.SUBCKT D1PS89SB74 1 2 3
*
* The resistors do not reflect
* physical devices. Instead they
* improve modeling in the reverse
* mode of operation.
*
R1 1 3 1.409E+09
D1 1 3 D1PS89SB74
R2 3 2 1.409E+09
D2 3 2 D1PS89SB74
*
.MODEL D1PS89SB74 D
+(
+    IS = 2.775E-09
+    N = 1.021
+    BV = 77
+    IBV = 1.67E-07
+    RS = 27.73
+    CJO = 1.655E-12
+    VJ = 0.349
+    M = 0.3583
+    FC = 0.5
+    TT = 0
+    EG = 0.69
+    XTI = 2
+)
.ENDS
*