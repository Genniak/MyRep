*BZT52C24 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*24V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C24 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  23.37
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=31.2P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=650U RS=21 N=9.5)
.ENDS