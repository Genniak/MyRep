*SI6331DQ  MCE  5-27-97
*30V 6A 0.025ohm Triple Power MOSFET pkg:SMD28 (A:1,4,26)(B:6,9,21)(C:11,14,16)
.SUBCKT SI6331DQ 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  10.9M
RS  40  3  1.63M
RG  20  2  26.8
CGS  2  3  1.3N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  517P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=1 KP=67.9)
.MODEL DCGD D (CJO=517P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=23.2N N=1.5 RS=1.79M BV=30 CJO=1.17N VJ=0.8 M=0.42 TT=50N)
.MODEL DLIM D (IS=100U)
.ENDS 