*SUP70N06-14 Siliconix 17-Mar-95
*N-Channel DMOS Subcircuit Model
.SUBCKT SUP70N06-14 4 1 2 2
M1 3 1 2 2 NMOS W=4251000U L=0.5U
R1 4 3 RTEMP 5.5M
CGS 1 2 1414PF
CGD 1 6 2700PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=80N RS=2M RD=0 LD=0
+ NSUB=4E+15 VTO=4.26 UO=350 VMAX=200K ETA=0.3M XJ=100N THETA=360M
+ KAPPA=0.05 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0 IS=0 NFS=0.5E+10)
.MODEL DMIN D(CJO=2300P VJ=0.08 M=0.48 FC=0.5 IS=1E-20 TT=10N)
.MODEL DMAX D(CJO=900P VJ=0.06 M=0.9 FC=0.5 IS=1E-16 TT=10N)
.MODEL DBODY D(CJO=1550P VJ=0.4 M=0.36 FC=0.5 N=1 IS=1E-15
+ TT=14N BV=68)
.MODEL RTEMP R(TC1=7M TC2=20U)
.ENDS 