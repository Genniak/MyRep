*ZPY10 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*10V 1.3W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZPY10    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  9.436
.MODEL DF D (IS=6.53N RS=32.3M N=1.7 CJO=89.6P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.41M RS=1.2 N=5.4)
.ENDS