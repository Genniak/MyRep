*
.SUBCKT BAT854SW 1 2 3
*
* The Resistor R1 does not reflect
* a physical device. Instead it
* improves modeling in the reverse
* mode of operation.
*
R1 1 3 9.5E+07
D1 1 3 BAT854SW
R2 3 2 9.5E+07
D2 3 2 BAT854SW
*
.MODEL BAT854SW D
+(
+ IS = 8E-08
+ N = 1.012
+ BV = 45
+ IBV = 0.0001
+ RS = 0.8243
+ CJO = 2.515E-11
+ VJ = 0.4182
+ M = 0.4941
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*