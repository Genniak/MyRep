*SI9934DY  MCE  5-28-97
* jjt 4/4/2002: changed sign of VTO to match S-49532�Rev. E, 02-Feb-98 datasheet
*12V 5A 0.045ohm Power MOSFET pkg:SMD8A (A:8,2,1)(B:6,4,3)
.SUBCKT SI9934DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  20.4M
RS  40  3  2.12M
RG  20  2  30
CGS  2  3  1.15N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  1.28N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=25K THETA=80M ETA=2M VTO=-0.6 KP=183)
.MODEL DCGD D (CJO=1.28N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=20.8N N=1.5 RS=0 BV=12 CJO=1.11N VJ=0.8 M=0.42 TT=67N)
.MODEL DLIM D (IS=100U)
.ENDS 