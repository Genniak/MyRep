*
.SUBCKT D1PS70SB20 1 2
* The Resistor R1 does not reflect
* a physical device. Instead it
* improves modeling in the reverse
* mode of operation.
*
R1 1 2 4.018E+06
D1 1 2 D1PS70SB20
*
.MODEL D1PS70SB20 D
+(
+ IS = 4.291E-06
+ N = 1.002
+ BV = 44
+ IBV = 3.0E-05
+ RS = 0.3772
+ CJO = 7.8E-11
+ VJ = 0.4015
+ M = 0.508
+ FC = 0.1
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*