*1N5347B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*10V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5347B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  9.415
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=68.9P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=7.18M RS=0.6 N=6.8)
.ENDS