*DL5236B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*7.5V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5236B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  6.964
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=53.1P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=52U RS=1.8 N=3.2)
.ENDS