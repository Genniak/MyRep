*DL5254B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*27V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5254B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  26.44
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=32.6P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=104U RS=12.3 N=5.1)
.ENDS