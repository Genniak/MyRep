*SI6802DQ  MCE  5-27-97
*20V 3A 0.057ohm Reduced Qg Power MOSFET pkg:SMD8B 1,4,6
.SUBCKT SI6802DQ 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  26.1M
RS  40  3  2.43M
RG  20  2  45.5
CGS  2  3  510P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  555P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=41.7K THETA=80M ETA=2M VTO=0.6 KP=80)
.MODEL DCGD D (CJO=555P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=300N N=1.5 RS=21.2M BV=20 CJO=1.06N VJ=0.8 M=0.42 TT=52N)
.MODEL DLIM D (IS=100U)
.ENDS 