*
.SUBCKT BAT74 1 2
* The resistors do not reflect
* physical devices.  Instead they
* improve modeling in the reverse
* mode of operation.
R1 1 2 2.9E+07
D1 1 2 BAT74
*
.MODEL BAT74 D
+(
+ IS = 2.548E-07
+ N = 1.02
+ BV = 33
+ IBV = 1.251E-06
+ RS = 2.582
+ CJO = 9.92E-12
+ VJ = 0.317
+ M = 0.4411
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*