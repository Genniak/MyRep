*
.SUBCKT BAT721S 1 2 3
* The resistors do not reflect
* physical devices. Instead they
* improve modeling in the reverse
* mode of operation.
R1 1 3 5.9E+06
D1 1 3 BAT721S
R2 3 2 5.9E+06
D2 3 2 BAT721S
*
.MODEL BAT721S D
+(
+ IS = 1.009E-06
+ N = 1.017
+ BV = 44
+ IBV = 0.001611
+ RS = 0.6578
+ CJO = 3.76E-11
+ VJ = 0.274
+ M = 0.4381
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*