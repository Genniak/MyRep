*DL5243B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*13V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5243B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  12.46
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=51.5P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=29.2U RS=3.9 N=3.3)
.ENDS