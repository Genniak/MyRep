*Si6953DQ Siliconix 13-Oct-94
*P-Channel DMOS Subcircuit Model
.SUBCKT Si6953DQ 4 1 2 2
M1 3 1 2 2 PMOS W=283290U L=0.5U
R1 4 3 RTEMP 40M
CGS 1 2 132PF
CGD 1 6 450PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=50N RS=56M RD=0 LD=0 NFS=3E+12
+ NSUB=8.7E+16 UO=110 VMAX=0 ETA=800U XJ=500N THETA=200U
+ KAPPA=0.3 CGBO=0 TPG=-1 DELTA=0.1 CGSO=0 CGDO=0 IS=0)
.MODEL DMIN D(CJO=380P VJ=0.25 M=0.58 FC=0.5)
.MODEL DMAX D(CJO=180P VJ=0.75 M=0.4 FC=0.5 IS=0.5E-24)
.MODEL DBODY D(CJO=590P VJ=0.35 M=0.335 FC=0.5 N=1 IS=1E-10
+ TT=14N BV=30)
.MODEL RTEMP R(TC1=13M TC2=0)
.ENDS Si6953DQ