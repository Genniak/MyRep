*ZY6_8 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*6.8V 2W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZY6_8    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  6.236
.MODEL DF D (IS=10N RS=21M N=1.7 CJO=246P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=2.81M RS=0.6 N=5.4)
.ENDS