*ZY82 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*82V 2W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZY82     1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  80.92
.MODEL DF D (IS=10N RS=21M N=1.7 CJO=38.2P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=4.9M RS=30 N=27)
.ENDS