*1N5386B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*180V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5386B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  178
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=20.3P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.59M RS=129 N=58)
.ENDS