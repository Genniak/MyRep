*Si4431DY Siliconix 26-Sep-95
*P-Channel DMOS Subcircuit Model
.SUBCKT Si4431DY 4 1 2 2
M1 3 1 2 2 PMOS W=1673620U L=0.5U
R1 4 3 RTEMP 10M
CGS 1 2 630PF
CGD 1 6 650PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=5E-8 RS=11M RD=0 LD=0 NFS=1.25E+12
+ NSUB=7.2E+16 UO=200 VMAX=0 ETA=1E-3 XJ=5E-7
+ KAPPA=1.5E-2 CGBO=0 THETA=0.5E-3 TPG=-1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=.065E-4)
.MODEL DMIN D(CJO=660E-12 VJ=0.25 M=0.4 FC=0.5)
.MODEL DMAX D(CJO=1080E-12 VJ=0.75 M=0.4 FC=0.5 IS=0.5E-15)
.MODEL DBODY D(CJO=1000E-12 VJ=0.35 M=0.335 FC=0.5 N=1 IS=5E-10
+ TT=6.0E-8 BV=40)
.MODEL RTEMP R(TC1=10E-3 TC2=1E-5)
.ENDS Si4431DY