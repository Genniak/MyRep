*DL5238B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*8.7V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5238B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  8.151
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=42.5P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=230U RS=2.4 N=4.3)
.ENDS