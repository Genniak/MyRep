*SI4946EY  MCE  5-27-97
*60V 4A 0.05ohm Dual Power MOSFET pkg:SMD8A (A:8,2,1)(B:6,4,3)
.SUBCKT SI4946EY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  22.8M
RS  40  3  2.25M
RG  20  2  33.3
CGS  2  3  880P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  327P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=125K THETA=80M ETA=2M VTO=1 KP=52.2)
.MODEL DCGD D (CJO=327P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=18.7N N=1.5 RS=33.3M BV=60 CJO=449P VJ=0.8 M=0.42 TT=35N)
.MODEL DLIM D (IS=100U)
.ENDS 