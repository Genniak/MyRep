*SI4450DY  MCE  5-27-97
*60V 8A 0.022ohm Power MOSFET pkg:SMD8A 8,4,1
.SUBCKT SI4450DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  9.45M
RS  40  3  1.55M
RG  20  2  20
CGS  2  3  1.54N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  725P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=125K THETA=80M ETA=2M VTO=2 KP=63.5)
.MODEL DCGD D (CJO=725P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=31.1N N=1.5 RS=0 BV=60 CJO=1.11N VJ=0.8 M=0.42 TT=46N)
.MODEL DLIM D (IS=100U)
.ENDS 