*
.SUBCKT BAS40-05W 1 2 3
* The Resistors do not
* reflect physical devices.
* Instead they improve modeling
* in the reverse mode of
* operation.
R1 1 3 6.659E+08
D1 1 3 BAS40-05W
R2 2 3 6.659E+08
D2 2 3 BAS40-05W
*
.MODEL BAS40-05W D
+(
+ IS = 1.419E-08
+ N = 1.025
+ BV = 44
+ IBV = 1.255E-07
+ RS = 4.942
+ CJO = 4.046E-12
+ VJ = 0.323
+ M = 0.4154
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*