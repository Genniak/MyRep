*Si4953DY Siliconix 13-Feb-96
*P-Channel DMOS Subcircuit Model
.SUBCKT Si4953DY 4 1 2 2
M1 3 1 2 2 PMOS W=1232400U L=0.5U
R1 4 3 RTEMP 21M
CGS 1 2 560PF
CGD 1 6 650PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=50N RS=20M RD=0 LD=0 NFS=0.8E+12
+ NSUB=7.4E+16 UO=200 VMAX=0 ETA=300U XJ=500N
+ KAPPA=0.1 CGBO=0 THETA=0 TPG=-1 DELTA=0 CGSO=0 CGDO=0
+ IS=0 KP=6.7U)
.MODEL DMIN D(CJO=560P VJ=0.22 M=0.42 FC=0.5 IS=1.0E-15)
.MODEL DMAX D(CJO=200P VJ=0.8 M=0.5 FC=0.5 IS=0.5E-15)
.MODEL DBODY D(CJO=790P VJ=0.7 M=0.4 FC=0.5 N=1 IS=1E-15
+ TT=1E-7 BV=40)
.MODEL RTEMP R(TC1=7.7M TC2=10U)
.ENDS Si4953DY