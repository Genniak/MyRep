*1N5345B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*8.7V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5345B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  8.092
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=85P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=13.9M RS=0.6 N=8.1)
.ENDS