*DL4751A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*30V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4751A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  29.37
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=46.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.04M RS=12 N=9.2)
.ENDS