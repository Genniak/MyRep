*
.SUBCKT BAT720 1 2
R1 1 2 2.8E+06
D1 1 2 DBAT720
*
* The Resistor R1 does not reflect
* a physical device.  Instead it
* improves modeling in the reverse
* mode of operation
*
.MODEL DBAT720 D
+(
+ IS = 1.281E-06
+ N = 1.009
+ BV = 44
+ IBV = 2.21E-05
+ RS = 0.3093
+ CJO = 8.133E-11
+ VJ = 0.4519
+ M = 0.5304
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*