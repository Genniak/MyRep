*Si4947DY Siliconix 01-Mar-96
*P-Channel DMOS Subcircuit Model
.SUBCKT Si4947DY 4 1 2 2
M1 3 1 2 2 PMOS W=648284U L=0.5U
R1 4 3 RTEMP 26M
CGS 1 2 270PF
CGD 1 6 400PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=5E-8 RS=30M RD=0 LD=0 NFS=1.25E+12
+ NSUB=7.2E+16 UO=200 VMAX=0 ETA=0.1M XJ=5E-7
+ KAPPA=9E-2 CGBO=0 THETA=1M TPG=-1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=6.15U)
.MODEL DMIN D(CJO=260P VJ=0.2 M=0.4 FC=0.5)
.MODEL DMAX D(CJO=180P VJ=0.75 M=0.4 FC=0.5 IS=0.5E-20)
.MODEL DBODY D(CJO=350P VJ=0.85 M=0.32 FC=0.5 N=1 IS=5E-14
+ TT=14.7E-8 BV=40)
.MODEL RTEMP R(TC1=12M TC2=25U)
.ENDS Si4947DY