*
.SUBCKT BAT721A 1 2 3
* The resistors do not reflect
* physical devices. Instead they
* improve modeling in the reverse
* mode of operation.
R1 3 1 5.9E+06
D1 3 1 BAT721A
R2 3 2 5.9E+06
D2 3 2 BAT721A
*
.MODEL BAT721A D
+(
+ IS = 1.009E-06
+ N = 1.017
+ BV = 44
+ IBV = 0.001611
+ RS = 0.6578
+ CJO = 3.76E-11
+ VJ = 0.274
+ M = 0.4381
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*