*
.SUBCKT D1PS76SBD17 1 2
* The Resistor R1 does not reflect
* a physical device.  Instead it
* improves modeling in the reverse
* mode of operation.
R1 1 2 6E+07
D1 1 2 SBD
.MODEL SBD D
+(
+ IS = 1.419E-09
+ N = 1.022
+ BV = 6
+ IBV = 2.45E-06
+ RS = 5.112
+ CJO = 7.867E-13
+ VJ = 0.1043
+ M = 0.1439
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*
*