*DL4746A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*18V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4746A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  17.4
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=67.8P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.09M RS=6 N=7.6)
.ENDS