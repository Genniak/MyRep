*SI9925DY  MCE  5-27-97
*20V 5A 0.045ohm Dual Power MOSFET pkg:SMD8A (A:8,2,1)(B:6,4,3)
.SUBCKT SI9925DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  20.4M
RS  40  3  2.12M
RG  20  2  30
CGS  2  3  720P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  634P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=41.7K THETA=80M ETA=2M VTO=0.8 KP=97.5)
.MODEL DCGD D (CJO=634P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=20.8N N=1.5 RS=12M BV=20 CJO=737P VJ=0.8 M=0.42 TT=60N)
.MODEL DLIM D (IS=100U)
.ENDS 