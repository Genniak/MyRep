*SI9426DY  MCE  5-27-97
*20V 10A 0.01ohm Power MOSFET pkg:SMD8A 1,4,6
.SUBCKT SI9426DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  3.75M
RS  40  3  1.25M
RG  20  2  15
CGS  2  3  2.86N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  179P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=41.7K THETA=80M ETA=2M VTO=0.6 KP=808)
.MODEL DCGD D (CJO=179P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=722N N=1.5 RS=7.1M BV=20 CJO=3.11N VJ=0.8 M=0.42 TT=59N)
.MODEL DLIM D (IS=100U)
.ENDS 