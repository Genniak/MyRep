*
.SUBCKT BAT721 1 3
* The resistor R1 does not reflect
* a physical device. Instead it
* improves modeling in the reverse
* mode of operation.
R1 1 3 5.9E+06
D1 1 3 BAT721
*
.MODEL BAT721 D
+(
+ IS = 1.009E-06
+ N = 1.017
+ BV = 44
+ IBV = 0.001611
+ RS = 0.6578
+ CJO = 3.76E-11
+ VJ = 0.274
+ M = 0.4381
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*