*ZY4_3 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*4.3V 2W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZY4_3    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  3.439
.MODEL DF D (IS=10N RS=21M N=1.7 CJO=489P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=36M RS=2.1 N=19)
.ENDS