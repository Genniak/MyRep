*DL5249B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*19V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5249B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  18.45
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=40P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=59.7U RS=6.9 N=4.1)
.ENDS