*ZPY16 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*16V 1.3W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZPY16    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  15.42
.MODEL DF D (IS=6.53N RS=32.3M N=1.7 CJO=92.2P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.44M RS=3 N=6.8)
.ENDS