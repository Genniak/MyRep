*
.SUBCKT D1PS75SB45 1 2 3
*
* The resistors do not reflect
* physical devices.  Instead they
* improve modeling in the reverse
* mode of operation.
*
R1 1 3 8E+08
D1 1 3 D1PS75SB45
R2 2 3 8E+08
D2 2 3 D1PS75SB45
.MODEL D1PS75SB45 D
+(
+ IS = 9.114E-09
+ N = 1.006
+ BV = 45
+ IBV = 7.8E-05
+ RS = 4.563
+ CJO = 3.895E-12
+ VJ = 0.3192
+ M = 0.4008
+ FC = 0.5
+ TT = 0
+ EG = 0.69
+ XTI = 2
+)
.ENDS
*