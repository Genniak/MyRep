*Si6946DQ Siliconix 22-Oct-96
*N-Channel DMOS Subcircuit Model
.SUBCKT Si6946DQ 4 1 2 2
M1 3 1 2 2 NMOS W=298454U L=0.5U
R1 4 3 RTEMP 45M
CGS 1 2 180PF
CGD 1 6 1165PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=17.5N RS=550U RD=0 LD=0
+ NSUB=2.6E+17 UO=800 VMAX=1MEG ETA=300U XJ=500N
+ KAPPA=0.25 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=80U NFS=0.8E+12)
.MODEL DMIN D(CJO=932P VJ=0.06 M=0.6 FC=0.5 IS=1E-18)
.MODEL DMAX D(CJO=860P VJ=0.6 M=0.5 FC=0.5 IS=1E-19)
.MODEL DBODY D(CJO=430P VJ=0.15 M=0.26 FC=0.5 N=1 IS=1E-15
+ TT=14N BV=40)
.MODEL RTEMP R(TC1=3.2M TC2=12U)
.ENDS 