*1N5380B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*120V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5380B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  118.4
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=22.9P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=6.57M RS=51 N=46)
.ENDS