*SUP65P06-20 Siliconix 01-May-95
*P-Channel DMOS Subcircuit Model
.SUBCKT SUP65P06-20 4 1 2 2
M1 3 1 2 2 PMOS W=4010100U L=0.5U
R1 4 3 RTEMP 6.7M
CGS 1 2 3410PF
CGD 1 6 2550PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=70N RS=4.2M RD=0 LD=0 NFS=1.1E+12
+ NSUB=1.25E+17 VTO=-1 UO=300 VMAX=0 ETA=100U XJ=1.7U THETA=1U
+ KAPPA=150M CGBO=0 TPG=-1 DELTA=0.1 CGSO=0 CGDO=0 IS=0)
.MODEL DMIN D(CJO=4180P VJ=0.15 M=0.5 FC=0.5)
.MODEL DMAX D(CJO=3000P VJ=0.95 M=0.4 FC=0.5 IS=0.5E-24)
.MODEL DBODY D(CJO=2450P VJ=0.5 M=0.38 FC=0.5 N=1 IS=1E-10
+ TT=14N BV=70)
.MODEL RTEMP R(TC1=9.5M TC2=5U)
.ENDS SUP65P06-20