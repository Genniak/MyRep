*Si9434DY Siliconix 21-Oct-96
*P-Channel DMOS Subcircuit Model
.SUBCKT Si9434DY 4 1 2 2
M1 3 1 2 2 PMOS W=1173406U L=0.5U
R1 4 3 RTEMP 10M
CGS 1 2 407PF
CGD 1 6 4231PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=17.5N RS=6M RD=0 LD=0
+ NSUB=4.86E+16 VTO=-1.38 UO=250 VMAX=0 ETA=300U XJ=500N THETA=0
+ KAPPA=5M CGBO=0 TPG=-1 DELTA=0 CGSO=0 CGDO=0 IS=0 KP=12.4U)
.MODEL DMIN D(CJO=4340P VJ=0.22 M=0.83 FC=0.56 IS=1E-20)
.MODEL DMAX D(CJO=1500P VJ=0.4 M=0.8 FC=0.5 IS=1E-22)
.MODEL DBODY D(CJO=1433P VJ=0.85 M=0.38 FC=0.5 N=1 IS=1E-18
+ TT=100N BV=20)
.MODEL RTEMP R(TC1=90M TC2=47U)
.ENDS Si9434DY