*Si6447DQ Siliconix 15-Nov-94
*P-Channel DMOS Subcircuit Model
.SUBCKT Si6447DQ 4 1 2 2
M1 3 1 2 2 PMOS W=492336U L=0.5U
R1 4 3 RTEMP 28M
CGS 1 2 146PF
CGD 1 6 950PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=30N RS=22M RD=0 LD=0 NFS=3E+12
+ NSUB=1.6E+17 UO=200 VMAX=0 ETA=0.8M XJ=500N
+ KAPPA=1E-1 CGBO=0 THETA=1U TPG=-1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=10.15U)
.MODEL DMIN D(CJO=880P VJ=0.25 M=0.58 FC=0.5)
.MODEL DMAX D(CJO=480P VJ=0.75 M=0.4 FC=0.5 IS=0.5E-24)
.MODEL DBODY D(CJO=990P VJ=0.35 M=0.335 FC=0.5 N=1 IS=1E-10
+ TT=14N BV=30)
.MODEL RTEMP R(TC1=10M TC2=0)
.ENDS Si6447DQ