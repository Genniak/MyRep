*SI4420DY  MCE  5-27-97
*30V 12A 0.0088ohm Power MOSFET pkg:SMD8A 8,4,1
.SUBCKT SI4420DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  3.18M
RS  40  3  1.22M
RG  20  2  12
CGS  2  3  4.6N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  4.13N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=1 KP=388)
.MODEL DCGD D (CJO=4.13N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=51.9N N=1.5 RS=20M BV=30 CJO=1.51N VJ=0.8 M=0.42 TT=49N)
.MODEL DLIM D (IS=100U)
.ENDS 