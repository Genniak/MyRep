*ZPY1 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*1V 1.3W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZPY1     1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  0.4881
.MODEL DF D (IS=6.53N RS=32.3M N=1.7 CJO=2.83N VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=87.8P RS=2.4 N=1.1)
.ENDS